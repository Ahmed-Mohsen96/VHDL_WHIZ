entity first_program is
-- define i/o 
end first_program;


architecture sim_f_program of first_program is
begin	
	process is
	begin
		report "Hello World !";
		wait;
	end process;



end sim_f_program;